
interface hbus_if;
	logic [`DATA-1:0] hdata;
	logic [`ADDR-1:0] addr;
	logic hen;
	logic hwr_rd;
endinterface
