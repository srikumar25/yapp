
package yapp_pkg;

`include "uvm_macros.svh"
import uvm_pkg::*;
`include "yapp_seq_item.sv"
`include "yapp_seq.sv"
`include "yapp_driver.sv"
`include "yapp_sequencer.sv"
//`include "yapp_monitor.sv"
//`include "yapp_agent_cfg.sv"
`include "yapp_agent.sv"
`include "yapp_env.sv"
//`include "yapp_test.sv"
`include "../test/yapp_basic_test.sv"

endpackage
