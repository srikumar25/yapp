
interface yapp_if;
	logic [`DATA-1:0] in_data;
	logic in_data_vld;
	logic in_suspend;
endinterface
