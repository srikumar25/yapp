
`ifndef YAPP_PKG
`define YAPP_PKG

//`include "../hbus/hbus_pkg.sv"
//`include "../chan/chan_pkg.sv"

package yapp_pkg;

`include "uvm_macros.svh"
import uvm_pkg::*;
import hbus_pkg::*;
import chan_pkg::*;
`include "yapp_seq_item.sv"
`include "yapp_driver.sv"
`include "yapp_sequencer.sv"
`include "yapp_agent_cfg.sv"
`include "yapp_agent.sv"
`include "yapp_monitor.sv"
//`include "yapp_test.sv"
`include "yapp_env.sv"
`include "../seq/hbus_basic_seq.sv"
`include "../../seq/yapp_basic_seq.sv"
`include "../../test/yapp_basic_test.sv"

endpackage
`endif
