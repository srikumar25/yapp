
interface chan_if;
	logic [`DATA-1:0] data;
	logic data_vld;
	logic suspend;
endinterface
