interface common;
	logic clk;
	logic rst;
	logic error;
endinterface
