
typedef uvm_sequencer#(yapp_seq_item) yapp_sequencer;
//typedef yapp_sequencer extends uvm_sequencer#(yapp_seq_item); 
//yapp_sequencer;

/*class yapp_sequencer extends uvm_sequencer;
	
	`uvm_component_utils(yapp_sequencer)

function void new("yapp_sequencer",null);
	super.new(yapp_sequencer,null);
endfunction

function void build_phase(uvm_phase phase);
	super.build_phase(phase);
endfunction

function void connect_phase(uvm_phase phase);
	super.connect_phase(phase);
endfunction

endclass 
*/
